module LM96570Control_NEW();

endmodule
