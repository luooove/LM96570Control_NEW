module LM96570(clk,reset_N,sRD,sLE,sWR,sCLK,TX_EN,RST);

//-------------与FPGA内部连接-------//
input clk; //时钟输入
input reset_N;// 复位信号


//-------------与硬件接口-------//
output sRD;  // 4-Wire Serial Interface Data Output for reading data registers
output sLE;  // 4-Wire Serial Interface Latch Enable
output sWR;  // 4-Wire Serial Interface Data Input for writing data registers
output sCLK; // 4-Wire Serial Interface Clock
output RST;  // Asynchronous Chip Reset
output TX_EN;//Beamformer starts firing

//-------------寄存器初始化-------//
reg addr_data; // 发送移位寄存其选择，1选地址移位寄存器，0选数据移位寄存器
reg [5:0]addr_buf; // 发送地址寄存器 5bits
reg [63:0]data_buf; // 发送数据寄存器 最大64bits

reg [4:0]addr_cfg[17:1]; // 具体地址member
reg [63:0]data_cfg[17:1]; // 具体数据member

//-------------计数器初始化-------//
reg [4:0]cnt_cfg;  // 配置计数器 输出几组数据（地址加数据）
reg [2:0]cnt_addr; // 地址位宽计数器
reg [5:0]cnt_data; // 数据位宽计数器

//-------------组合逻辑处理-------//
assign sWR  = addr_data?addr_buf[0]:data_buf[0]; //1选地址移位寄存器，0选数据移位寄存器
assign sCLK = link_sCLK?clk:1'b0; 

//-------------状态机初始化-------//
reg state[5:0];
parameter   IDLE        = 6'000_001;
				ADDR_OUT		= 6'000_010; 
				DATA_OUT		= 6'000_100; 
				DATA_IN		= 6'001_000; 
				ACK_OUT		= 6'010_000; 
				ACK_IN		= 6'100_000; 

//-------------开关定义-------//
parameter YES  =1'b1,
          NO   =1'b0;

			 
			 
//------------主状态机程序-------//
always@(negedge clk or negedge reset_N)
if(!reset_N) //系统复位初始化
	begin
		addr_cfg[17]<=5'b11010;            //地址1A
		//addr_cfg[2]<=5'b11001;            //地址19
		//addr_cfg[1]<=5'b11000;            //地址18
		

		addr_cfg[16]<=5'b10111;            //地址17h
		addr_cfg[15]<=5'b10111;            //地址16h
		addr_cfg[14]<=5'b10111;            //地址15h
		addr_cfg[13]<=5'b10111;            //地址14h
		addr_cfg[12]<=5'b10111;            //地址13h
		addr_cfg[11]<=5'b10111;            //地址12h
		addr_cfg[10]<=5'b10111;            //地址11h
		addr_cfg[9]<=5'b10111;            //地址10h
		
		addr_cfg[8]<=5'b10111;            //地址0Fh
		addr_cfg[7]<=5'b10111;            //地址0Eh
		addr_cfg[6]<=5'b10111;            //地址0Dh
		addr_cfg[5]<=5'b10111;            //地址0Ch
		addr_cfg[4]<=5'b10111;            //地址0Bh
		addr_cfg[3]<=5'b10111;            //地址0Ah
		addr_cfg[2]<=5'b10111;            //地址09h
		addr_cfg[1]<=5'b01111;            //地址08h
		
		data_cfg[17]<=64'b0000_0000_0000_0000__0000_0000_0000_0000__0000_0000_0000_000000__00_0110_0000_0111;
		//data_cfg[2]<=64'b1111_0000_1111_1110__0000_0011_1111_0000__0011_1110_0000_1111__0000_1110_0011_0010;
		//data_cfg[1]<=64'b0000_1111_0000_0001__1111_1100_0000_1111__1100_0001_1111_0000__1111_0001_1100_1101;
		data_cfg[16]<=64'b0000_0000_0000_0000__0000_0000_0000_0000__0000_0000_0000_0000__0000_0000_0000_0000;
		data_cfg[15]<=64'b0000_0000_0000_0000__0000_0000_0000_0000__0000_0000_0000_0000__0000_0000_0000_0000;
		data_cfg[14]<=64'b0000_0000_0000_0000__0000_0000_0000_0000__0000_0000_0000_0000__0000_0000_0000_0000;
		data_cfg[13]<=64'b0000_0000_0000_0000__0000_0000_0000_0000__0000_0000_0000_0000__0000_0000_0000_0000;
		data_cfg[12]<=64'b0000_0000_0000_0000__0000_0000_0000_0000__0000_0000_0000_0000__0000_0000_0000_0000;
		data_cfg[11]<=64'b0000_0000_0000_0000__0000_0000_0000_0000__0000_0000_0000_0000__0000_0000_0000_0000;
		data_cfg[10]<=64'b0000_0000_0000_0000__0000_0000_0000_0000__0000_0000_0000_0000__0000_0000_0000_0000;
		data_cfg[9]<=64'b0101_0101_0101_0101__0101_0101_0101_0101__0101_0101_0101_0101__0101_0101_0101_0101;
		data_cfg[8]<=64'b0000_0000_0000_0000__0000_0000_0000_0000__0000_0000_0000_0000__0000_0000_0000_0000;
		data_cfg[7]<=64'b0000_0000_0000_0000__0000_0000_0000_0000__0000_0000_0000_0000__0000_0000_0000_0000;
		data_cfg[6]<=64'b0000_0000_0000_0000__0000_0000_0000_0000__0000_0000_0000_0000__0000_0000_0000_0000;
		data_cfg[5]<=64'b0000_0000_0000_0000__0000_0000_0000_0000__0000_0000_0000_0000__0000_0000_0000_0000;
		data_cfg[4]<=64'b0000_0000_0000_0000__0000_0000_0000_0000__0000_0000_0000_0000__0000_0000_0000_0000;
		data_cfg[3]<=64'b0000_0000_0000_0000__0000_0000_0000_0000__0000_0000_0000_0000__0000_0000_0000_0000;
		data_cfg[2]<=64'b0000_0000_0000_0000__0000_0000_0000_0000__0000_0000_0000_0000__0000_0000_0000_0000;
		//data_cfg[1]<=64'b0101_0101_0101_0101__0101_0101_0101_0101__0101_0101_0101_0101__0101_0101_0101_0101;
		data_cfg[1]<=64'b1010_1010_1010_1010__1010_1010_1010_1010__1010_1010_1010_1010__1010_1010_1010_1010;
		
		TX_EN	   <= NO;
		sLE      <= 1'b1;
		cnt_cfg  <= 5'b1001; //17
		state    <= IDLE;
		
	end
else	
	begin
		casex(state)
			IDLE:begin
						sLE <= 1'b1;
						link sCLK <= NO;
						link_sWR <= NO;
						addr_data <= 1'b1; //输出地址
						if(cnt_cfg)
							begin
								addr_buf <= {1'b0,addr_cfg[cnt_cfg]};
								data_buf <= data_cfg[cnt_cfg];
								TX_EN 	<= NO;
								state		<= ADDR_OUT;
							end
					end
			ADDR_OUT:begin
						sLE 		 <= 1'b0;
						link_sCLK <= YES;
						link_sWR	 <= YES;
						cnt_addr  <=3'b101;  //5
						casex(addr_buf[4:0])   //不同的地址位宽不一样，进行判断
							5'b00???:cnt_data<=6'b01_0101;  //21
							5'b01???:cnt_data<=6'b11_1111;  //63
							5'b10???:cnt_data<=6'b11_1111;  //63
							5'b1100?:cnt_data<=6'b11_1111;  //63
							5'b11010:cnt_data<=6'b00_1101;  //13
						endcase
						cnt_cfg<=cnt_cfg-1'b1;
						state<=DATA_OUT;
					end
			DATA_OUT:begin
							if(cnt_addr)
								begin
								   addr_buf<=addr_buf>>1'b1;
									cnt_addr<=cnt_addr-1'b1;
								end
					end
					
	end

	

				
endmodule
